`ifndef __SYS_DEFS_SVH__
`define __SYS_DEFS_SVH__
`timescale 1ns/1ps

`define DATA_LEN 31
`define MEMDEPTH 31
`define SHIFT_LEN 5
